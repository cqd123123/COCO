module DataExtension(input [31:0] Din,input [2:0] ExtFunct,input [1:0] A1_A0,output [31:0] ExtDout);
  assign ExtDout=(ExtFunct==3'b001)?
                ((A1_A0==2'b00)?{24'b00000000_00000000_00000000,Din[7:0]}:
                (A1_A0==2'b01)?{24'b00000000_00000000_00000000,Din[15:8]}:
                (A1_A0==2'b10)?{24'b00000000_00000000_00000000,Din[23:16]}:
                (A1_A0==2'b11)?{24'b00000000_00000000_00000000,Din[31:24]}:Din)
                :
                (ExtFunct==3'b010)?
                ((A1_A0==2'b00)?{16'b00000000_00000000,Din[15:0]}:
                (A1_A0==2'b10)?{16'b00000000_00000000,Din[31:16]}:Din)
                :
                (ExtFunct==3'b011)?
                ((A1_A0==2'b00)?{{24{Din[7]}},Din[7:0]}:
                (A1_A0==2'b01)?{{24{Din[15]}},Din[15:8]}:
                (A1_A0==2'b10)?{{24{Din[23]}},Din[23:16]}:
                (A1_A0==2'b11)?{{24{Din[31]}},Din[31:24]}:Din)
                :
                (ExtFunct==3'b100)?
                ((A1_A0==2'b00)?{{16{Din[15]}},Din[15:0]}:
                (A1_A0==2'b10)?{{16{Din[31]}},Din[31:16]}:Din)
                :Din;           
endmodule
