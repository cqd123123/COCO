module ALU(input [31:0] A,B,input [3:0] Ctrl,output [31:0] C,output Zero,Overflow,Compare);
  assign C=(Ctrl==4'b1110)?{B[15:0],16'h0000}://lui
           (Ctrl==4'b0000)?(A+B):
           (Ctrl==4'b0001)?(A+B)://
           (Ctrl==4'b0010)?(A-B):
           (Ctrl==4'b0011)?(A-B)://
           (Ctrl==4'b0100)?A&B:
           (Ctrl==4'b0101)?A|B:
           (Ctrl==4'b0110)?~(A|B)://nor
           (Ctrl==4'b0111)?A^B:
           (Ctrl==4'b1000)?((A<B)?1:0): //sltu
           (Ctrl==4'b1001)?   //slt
           (((A[31]==0&&B[31]==0)||(A[31]==1&&B[31]==1))?((A<B)?32'h00000001:32'h00000000):
           (A[31]==1&&B[31]==0)?32'h00000001:
           (A[31]==0&&B[31]==1)?32'h00000000:32'hffffffff)
           :32'hffffffff;
  assign Compare=(Ctrl==4'b1010)?((A[31]==1)?1:0):
                 (Ctrl==4'b1011)?(((A[31]==1)||(|A[31:0]==0))?1:0):
                 (Ctrl==4'b1100)?(((A[31]==0)&&(|A[31:0]!=0))?1:0):
                 (Ctrl==4'b1101)?((A[31]==0)?1:0):0;
  assign Zero=~(|C[31:0]);
  assign Overflow=(Ctrl==4'b0001)?(((A[31]==0&&B[31]==0&&C[31]==1)||(A[31]==1&&B[31]==1&&C[31]==0))?1:0):
                  (Ctrl==4'b0011)?(((A[31]==0&&B[31]==1&&C[31]==1)||(A[31]==1&&B[31]==0&&C[31]==1))?1:0):0;
endmodule